LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY EX6 IS
	PORT(CLK,CLR:IN STD_LOGIC;OPT:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END ENTITY EX6;

ARCHITECTURE LOGIC OF EX6 IS
SIGNAL CURRENT_DATA:STD_LOGIC_VECTOR(3 DOWNTO 0):="0000";
BEGIN

	PROCESS(CLK,CLR)
	BEGIN
		IF(CLR='1')THEN
			CURRENT_DATA<="0000";
		ELSIF(CLK'EVENT AND CLK='1')THEN
			IF (CURRENT_DATA="1001")THEN
				CURRENT_DATA<="0000";
			ELSE
				CURRENT_DATA<=CURRENT_DATA+1;
			END IF;
		END IF;
	END PROCESS;
	
	OPT <= "1111110" WHEN CURRENT_DATA = "0000" ELSE
		"0110000" WHEN CURRENT_DATA = "0001" ELSE
		"1101101" WHEN CURRENT_DATA = "0010" ELSE
		"1111001" WHEN CURRENT_DATA = "0011" ELSE
		"0110011" WHEN CURRENT_DATA = "0100" ELSE
		"1011011" WHEN CURRENT_DATA = "0101" ELSE
		"1011111" WHEN CURRENT_DATA = "0110" ELSE
		"1110000" WHEN CURRENT_DATA = "0111" ELSE
		"1111111" WHEN CURRENT_DATA = "1000" ELSE
		"1111011" WHEN CURRENT_DATA = "1001";
	
END LOGIC;